
`ifndef __RSTGEN_SEQUENCER_SV__
`define __RSTGEN_SEQUENCER_SV__

`include "rstgen_sequencer.svh"

function void rstgen_sequencer::build_phase(uvm_phase phase);
    super.build_phase(phase);
endfunction: build_phase

`endif //__RSTGEN_SEQUENCER_SV__
