
`ifndef __RSTGEN_PKG_SV__
`define __RSTGEN_PKG_SV__

`timescale 1ns / 1ps

package rstgen_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "rstgen_config.sv"
    `include "rstgen_transaction.sv"
    `include "rstgen_sequencer.sv"
    `include "rstgen_sequence.sv"
    `include "rstgen_monitor.sv"
    `include "rstgen_driver.sv"
    `include "rstgen_agent.sv"

endpackage: rstgen_pkg
`endif //__RSTGEN_PKG_SV__
